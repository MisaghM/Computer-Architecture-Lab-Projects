module RegsIdEx();

endmodule
