module StageId(
    input clk, rst,
    input [31:0] pcIn,
    output [31:0] pcOut
);
    assign pcOut = pcIn;
endmodule
