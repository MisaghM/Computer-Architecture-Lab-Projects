module InstructionDecode();

endmodule
