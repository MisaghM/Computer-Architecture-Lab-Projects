module RegsMemWb();

endmodule
