module Execution();

endmodule
