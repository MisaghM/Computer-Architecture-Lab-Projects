module WriteBack();

endmodule
