module RegsIfId();

endmodule
