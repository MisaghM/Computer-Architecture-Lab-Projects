module RegsExMem();

endmodule
