module RegsIfId(
    input clk, rst,
    input freeze, flush,
    input [31:0] pcIn, instructionIn,
    output reg [31:0] pcOut, instructionOut
);

endmodule
