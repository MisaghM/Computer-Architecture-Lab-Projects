module Memory();

endmodule
